module coefficients
(
	input logic [4:0] i_idx,
	output logic [15:0] o_tap
);

logic [3:0] state, next_state; // counter for which coefficient to send
logic [15:0] [15:0] taps; // array for 16 taps, just for testing

initial begin // initialize taps array for sim
	taps = '{'{1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1},
			'{1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1},
			'{1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1},
			'{1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1},
			'{1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1},
			'{1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1},
			'{1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1},
			'{1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1},
			'{1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1},
			'{1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1},
			'{1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1},
			'{1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1},
			'{1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1},
			'{1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1},
			'{1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1},
			'{1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1}};
end

always_comb begin
	o_tap = taps[15:0][i_idx];
end

endmodule